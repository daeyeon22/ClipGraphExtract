###############################################################################
#TSMC Library/IP Product
#Filename: tcbn65gplus_m8T2.lef
#Technology: CLN65GPLUS
#Product Type: Standard Cell
#Product Name: tcbn65gplus
#Version: 120a
###############################################################################
# 
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
# 
###############################################################################

# Resistor & Capacitor are referenced from spice model interconnect table
# The index is "width=minWidth", "Space=Pitch"
VERSION	5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
    CAPACITANCE PICOFARADS 10 ;
    CURRENT MILLIAMPS 10000 ;
    VOLTAGE VOLTS 1000 ;
    FREQUENCY MEGAHERTZ 10 ;
    DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER PO
    TYPE MASTERSLICE ;
END PO

LAYER CO
    TYPE CUT ;
END CO

PROPERTYDEFINITIONS 
    LAYER LEF57_SPACING STRING ;
END PROPERTYDEFINITIONS 

LAYER M1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.200 ;
    OFFSET 0.000 ;
    HEIGHT 0.5900 ;
    THICKNESS 0.1800 ;
    MINSTEP 0.090 ; 
    FILLACTIVESPACING 0.300 ;
    WIDTH 0.09 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    0.38    0.42    1.50    4.50
    WIDTH    0.00         0.09    0.09    0.09    0.09    0.09
    WIDTH    0.20         0.09    0.11    0.11    0.11    0.11
    WIDTH    0.42         0.09    0.11    0.16    0.16    0.16
    WIDTH    1.50         0.09    0.11    0.16    0.50    0.50
    WIDTH    4.50         0.09    0.11    0.16    0.50    1.50 ;
    PROPERTY LEF57_SPACING "SPACING 0.11 ENDOFLINE 0.11 WITHIN 0.035 PARALLELEDGE 0.11 WITHIN 0.11 ;" ;
    AREA 0.042 ;
    MINENCLOSEDAREA 0.20 ;

    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;
 
    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;

    MINIMUMCUT 2 WIDTH 0.300 ;
    MINIMUMCUT 4 WIDTH 0.700 ;
    MINIMUMCUT 2 WIDTH 0.300 LENGTH 0.300 WITHIN 0.800 ;
    MINIMUMCUT 2 WIDTH 2.000 LENGTH 2.000 WITHIN 2.000 ;
    MINIMUMCUT 2 WIDTH 3.000 LENGTH 10.000 WITHIN 5.000 ;

    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;

    ACCURRENTDENSITY 	AVERAGE
        FREQUENCY 	500 ;
        WIDTH     	0.090 	1.000 ;
        TABLEENTRIES	1.241	1.485 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH		0.090	0.180	0.500	1.000	5.000	12.000 ;
        TABLEENTRIES	14.936	13.727	11.656	10.736	9.829	9.681 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.090 1.0 12 ;
        TABLEENTRIES	41.861 50.097 50.844 ;
    RESISTANCE RPERSQ 0.1600000000 ;
    CAPACITANCE CPERSQDIST 0.0001711111 ;
    EDGECAPACITANCE 0.0000883000 ;
END M1

LAYER VIA1
    TYPE CUT ;
    SPACING 0.10 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    PROPERTY LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
    ANTENNAAREARATIO        20.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	15.8 ;
END VIA1

LAYER M2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.200 ;
    OFFSET 0.100 ;
    HEIGHT 0.9450 ;
    THICKNESS 0.2200 ;
    MINSTEP 0.100 ;
    FILLACTIVESPACING 0.300 ;
    WIDTH 0.1 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    0.38    0.40    1.50    4.50
    WIDTH    0.00         0.10    0.10    0.10    0.10    0.10
    WIDTH    0.20         0.10    0.12    0.12    0.12    0.12
    WIDTH    0.40         0.10    0.12    0.16    0.16    0.16
    WIDTH    1.50         0.10    0.12    0.16    0.50    0.50
    WIDTH    4.50         0.10    0.12    0.16    0.50    1.50 ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    AREA 0.052 ;
    MINENCLOSEDAREA 0.20 ;   

    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;
 
    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;

    MINIMUMCUT 2 WIDTH 0.300 ;
    MINIMUMCUT 4 WIDTH 0.700 ;
    MINIMUMCUT 2 WIDTH 0.300 LENGTH 0.300 WITHIN 0.800 ;
    MINIMUMCUT 2 WIDTH 2.000 LENGTH 2.000 WITHIN 2.000 ;
    MINIMUMCUT 2 WIDTH 3.000 LENGTH 10.000 WITHIN 5.000 ;

    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
  
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH		0.100	1.000 ;
        TABLEENTRIES 	1.577	1.847 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH     	0.100	0.200	0.500	1.000	5.000	12.000 ;
        TABLEENTRIES	9.324	8.384	7.101	6.451	5.803	5.696 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.100 1.0 12 ;
        TABLEENTRIES	26.135 30.615 31.071 ;
                		
    RESISTANCE RPERSQ 0.1400000000 ;
    CAPACITANCE CPERSQDIST 0.0002320000 ;
    EDGECAPACITANCE 0.0000780000 ;
END M2

LAYER VIA2
    TYPE CUT ;
    SPACING 0.10 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    PROPERTY LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
    ANTENNAAREARATIO        20.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	15.8 ;
END VIA2

LAYER M3
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.200 ;
    OFFSET 0.000 ;
    HEIGHT 1.3400 ;
    THICKNESS 0.2200 ;
    MINSTEP 0.100 ;
    FILLACTIVESPACING 0.300 ;
    WIDTH 0.1 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    0.38    0.40    1.50    4.50
    WIDTH    0.00         0.10    0.10    0.10    0.10    0.10
    WIDTH    0.20         0.10    0.12    0.12    0.12    0.12
    WIDTH    0.40         0.10    0.12    0.16    0.16    0.16
    WIDTH    1.50         0.10    0.12    0.16    0.50    0.50
    WIDTH    4.50         0.10    0.12    0.16    0.50    1.50 ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    AREA 0.052 ;
    MINENCLOSEDAREA 0.20 ;   

    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;
 
    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;

    MINIMUMCUT 2 WIDTH 0.300 ;
    MINIMUMCUT 4 WIDTH 0.700 ;
    MINIMUMCUT 2 WIDTH 0.300 LENGTH 0.300 WITHIN 0.800 ;
    MINIMUMCUT 2 WIDTH 2.000 LENGTH 2.000 WITHIN 2.000 ;
    MINIMUMCUT 2 WIDTH 3.000 LENGTH 10.000 WITHIN 5.000 ;

    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
  
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH		0.100	1.000 ;
        TABLEENTRIES 	1.577	1.847 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH     	0.100	0.200	0.500	1.000	5.000	12.000 ;
        TABLEENTRIES	8.965	7.789	6.191	5.347	4.453	4.299 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.100 1.0 12 ;
        TABLEENTRIES	26.135 30.615 31.071 ;
              		
    RESISTANCE RPERSQ 0.1400000000 ;
    CAPACITANCE CPERSQDIST 0.0002320000 ;
    EDGECAPACITANCE 0.0000779000 ;
END M3

LAYER VIA3
    TYPE CUT ;
    SPACING 0.10 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    PROPERTY LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
    ANTENNAAREARATIO        20.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	15.8 ;
END VIA3

LAYER M4
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.200 ;
    OFFSET 0.100 ;
    HEIGHT 1.7350 ;
    THICKNESS 0.2200 ;
    MINSTEP 0.100 ;
    FILLACTIVESPACING 0.300 ;
    WIDTH 0.1 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    0.38    0.40    1.50    4.50
    WIDTH    0.00         0.10    0.10    0.10    0.10    0.10
    WIDTH    0.20         0.10    0.12    0.12    0.12    0.12
    WIDTH    0.40         0.10    0.12    0.16    0.16    0.16
    WIDTH    1.50         0.10    0.12    0.16    0.50    0.50
    WIDTH    4.50         0.10    0.12    0.16    0.50    1.50 ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    AREA 0.052 ;
    MINENCLOSEDAREA 0.20 ;   

    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;
 
    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;
  
    MINIMUMCUT 2 WIDTH 0.300 ;
    MINIMUMCUT 4 WIDTH 0.700 ;
    MINIMUMCUT 2 WIDTH 0.300 LENGTH 0.300 WITHIN 0.800 ;
    MINIMUMCUT 2 WIDTH 2.000 LENGTH 2.000 WITHIN 2.000 ;
    MINIMUMCUT 2 WIDTH 3.000 LENGTH 10.000 WITHIN 5.000 ;
  
    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
  
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH		0.100	1.000 ;
        TABLEENTRIES 	1.577	1.847 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH     	0.100	0.200	0.500	1.000	5.000	12.000 ;
        TABLEENTRIES	8.824	7.548	5.805	4.857	3.811	3.623 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.100 1.0 12 ;
        TABLEENTRIES	26.135 30.615 31.071 ;

    RESISTANCE RPERSQ 0.1400000000 ;
    CAPACITANCE CPERSQDIST 0.0002320000 ;
    EDGECAPACITANCE 0.0000778000 ;
END M4

LAYER VIA4
    TYPE CUT ;
    SPACING 0.10 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    PROPERTY LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
    ANTENNAAREARATIO        20.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	15.8 ;
END VIA4

LAYER M5
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.200 ;
    OFFSET 0.000 ;
    HEIGHT 2.1300 ;
    THICKNESS 0.2200 ;
    MINSTEP 0.100 ;
    FILLACTIVESPACING 0.300 ;
    WIDTH 0.1 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    0.38    0.40    1.50    4.50
    WIDTH    0.00         0.10    0.10    0.10    0.10    0.10
    WIDTH    0.20         0.10    0.12    0.12    0.12    0.12
    WIDTH    0.40         0.10    0.12    0.16    0.16    0.16
    WIDTH    1.50         0.10    0.12    0.16    0.50    0.50
    WIDTH    4.50         0.10    0.12    0.16    0.50    1.50 ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    AREA 0.052 ;
    MINENCLOSEDAREA 0.20 ;   

    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;
 
    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;
  
    MINIMUMCUT 2 WIDTH 0.300 ;
    MINIMUMCUT 4 WIDTH 0.700 ;
    MINIMUMCUT 2 WIDTH 0.300 LENGTH 0.300 WITHIN 0.800 ;
    MINIMUMCUT 2 WIDTH 2.000 LENGTH 2.000 WITHIN 2.000 ;
    MINIMUMCUT 2 WIDTH 3.000 LENGTH 10.000 WITHIN 5.000 ;
  
    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
  
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH		0.100	1.000 ;
        TABLEENTRIES 	1.577	1.847 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH     	0.100	0.200	0.500	1.000	5.000	12.000 ;
        TABLEENTRIES	8.752	7.421	5.592	4.578	3.423	3.208 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.100 1.0 12 ;
        TABLEENTRIES	26.135 30.615 31.071 ;

    RESISTANCE RPERSQ 0.1400000000 ;
    CAPACITANCE CPERSQDIST 0.0002320000 ;
    EDGECAPACITANCE 0.0000778000 ;
END M5

LAYER VIA5
    TYPE CUT ;
    SPACING 0.10 ;
    SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
    PROPERTY LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
    ANTENNAAREARATIO        20.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	15.8 ;
END VIA5

LAYER M6
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.200 ;
    OFFSET 0.100 ;
    HEIGHT 2.5250 ;
    THICKNESS 0.2200 ;
    MINSTEP 0.100 ;
    FILLACTIVESPACING 0.300 ;
    WIDTH 0.1 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    0.38    0.40    1.50    4.50
    WIDTH    0.00         0.10    0.10    0.10    0.10    0.10
    WIDTH    0.20         0.10    0.12    0.12    0.12    0.12
    WIDTH    0.40         0.10    0.12    0.16    0.16    0.16
    WIDTH    1.50         0.10    0.12    0.16    0.50    0.50
    WIDTH    4.50         0.10    0.12    0.16    0.50    1.50 ;
    PROPERTY LEF57_SPACING "SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;" ;
    AREA 0.052 ;
    MINENCLOSEDAREA 0.20 ;   

    MINIMUMDENSITY 15 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 70 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;
 
    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;
  
    MINIMUMCUT 2 WIDTH 0.300 FROMBELOW ;
    MINIMUMCUT 4 WIDTH 0.700 FROMBELOW ;
    MINIMUMCUT 2 WIDTH 0.300 FROMBELOW LENGTH 0.300 WITHIN 0.800 ;
    MINIMUMCUT 2 WIDTH 2.000 FROMBELOW LENGTH 2.000 WITHIN 2.000 ;
    MINIMUMCUT 2 WIDTH 3.000 FROMBELOW LENGTH 10.000 WITHIN 5.000 ;
    MINIMUMCUT 2 WIDTH 1.800 FROMABOVE ;
    MINIMUMCUT 2 WIDTH 3.000 FROMABOVE LENGTH 10.0 WITHIN 5.001 ;
  
    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
  
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH		0.100   1.000 ;
        TABLEENTRIES 	1.577	1.847 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH     	0.100	0.200	0.500	1.000	5.000	12.000 ;
        TABLEENTRIES	8.701	7.336	5.453	4.394	3.158	2.921 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.100 1.0 12 ;
        TABLEENTRIES	26.135 30.615 31.071 ;

    RESISTANCE RPERSQ 0.1400000000 ;
    CAPACITANCE CPERSQDIST 0.0002320000 ;
    EDGECAPACITANCE 0.0000778000 ;
END M6

LAYER VIA6
    TYPE CUT ;
    SPACING 0.340 ;
    SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.56 ;
    ANTENNAAREARATIO        20.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	23.742 ;
END VIA6

LAYER M7
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.800 ;
    OFFSET 0.000 ;
    HEIGHT 3.3400 ;
    THICKNESS 0.9000 ;
    MINSTEP 0.400 ;
    FILLACTIVESPACING 0.600 ;
    WIDTH 0.400 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    1.50    4.50
    WIDTH    0.00         0.40    0.40    0.40
    WIDTH    1.50         0.40    0.50    0.50
    WIDTH    4.50         0.40    0.50    1.50 ;
    AREA 0.565 ;
    MINENCLOSEDAREA 0.565 ;   

    MINIMUMDENSITY 20 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 80 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;

    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;
  
    MINIMUMCUT 2 WIDTH 1.800 ;
    MINIMUMCUT 2 WIDTH 3.000 LENGTH 10.0 WITHIN 5.001 ;
  
    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 50480 ) ( 0.5 54000 ) ( 1 58000 ) ( 1.5 62000 ) ) ;
  
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH		0.400	1.000 ;
        TABLEENTRIES 	7.691	7.934 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH     	0.400	0.600	0.800	1.000	5.000	12.000 ;
        TABLEENTRIES	11.490	9.972	9.037	8.396	5.667	5.116 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.400 1.0 12 ;
        TABLEENTRIES	84.641 87.314 88.947 ;
  
    RESISTANCE RPERSQ 0.0220000000 ;
    CAPACITANCE CPERSQDIST 0.0000632500 ;
    EDGECAPACITANCE 0.0000915000 ;
END M7

LAYER VIA7
    TYPE CUT ;
    SPACING 0.340 ;
    SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.56 ;
    ANTENNAAREARATIO        20.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	23.742 ;
END VIA7

LAYER M8
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.800 ;
    OFFSET 0.100 ;
    HEIGHT 5.0400 ;
    THICKNESS 0.9000 ;
    MINSTEP 0.400 ;
    FILLACTIVESPACING 0.600 ;
    WIDTH 0.400 ;
    MAXWIDTH 12.0 ;
    SPACINGTABLE
    PARALLELRUNLENGTH     0.00    1.50    4.50
    WIDTH    0.00         0.40    0.40    0.40
    WIDTH    1.50         0.40    0.50    0.50
    WIDTH    4.50         0.40    0.50    1.50 ;
    AREA 0.565 ;
    MINENCLOSEDAREA 0.565 ;   

    MINIMUMDENSITY 20 ;
    MAXIMUMDENSITY 100 ;
    DENSITYCHECKWINDOW 50 50 ;
    DENSITYCHECKSTEP 25 ;
 
    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 80 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP 50 ;

    MINIMUMDENSITY 0 ;
    MAXIMUMDENSITY 90 ;
    DENSITYCHECKWINDOW 20 20 ;
    DENSITYCHECKSTEP 10 ;
  
    MINIMUMCUT 2 WIDTH 1.800 ;
    MINIMUMCUT 2 WIDTH 3.000 LENGTH 10.0 WITHIN 5.001 ;
  
    ANTENNACUMAREARATIO     5000.000000 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 50480 ) ( 0.5 54000 ) ( 1 58000 ) ( 1.5 62000 ) ) ;
  
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH		0.400	1.000 ;
        TABLEENTRIES 	7.691	7.934 ;
    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH     	0.400	0.600	0.800	1.000	5.000	12.000 ;
        TABLEENTRIES	11.373	9.827	8.870	8.213	5.372	4.783 ;
    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH		0.400 1.0 12 ;
        TABLEENTRIES	84.641 87.314 88.947 ;

    RESISTANCE RPERSQ 0.0220000000 ;
    CAPACITANCE CPERSQDIST 0.0000632500 ;
    EDGECAPACITANCE 0.0000956000 ;
END M8

LAYER OVERLAP
    TYPE OVERLAP ;
END OVERLAP

VIA VIA12_1cut DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M1 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA12_1cut

VIA VIA12_1cut_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M1 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA12_1cut_H
                 
VIA VIA12_1cut_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M1 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA12_1cut_V

VIA VIA12_1cut_FAT_C DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M1 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA12_1cut_FAT_C
             
VIA VIA12_1cut_FAT_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M1 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA12_1cut_FAT_H

VIA VIA12_1cut_FAT_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M1 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA12_1cut_FAT_V

VIA VIA12_1cut_FAT DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M1 ;
        RECT -0.090 -0.090  0.090  0.090 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M2 ;
        RECT -0.090 -0.090  0.090  0.090 ;
END VIA12_1cut_FAT
                 
VIA VIA12_2cut_E DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M1 ;
        RECT -0.090 -0.050  0.290  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.250  0.090 ;
END VIA12_2cut_E

VIA VIA12_2cut_W DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M1 ;
        RECT -0.290 -0.050  0.090  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M2 ;
        RECT -0.250 -0.090  0.050  0.090 ;
END VIA12_2cut_W

VIA VIA12_2cut_N DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M1 ;
        RECT -0.090 -0.050  0.090  0.250 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.290 ;
END VIA12_2cut_N

VIA VIA12_2cut_S DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M1 ;
        RECT -0.090 -0.250  0.090  0.050 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M2 ;
        RECT -0.050 -0.290  0.050  0.090 ;
END VIA12_2cut_S

VIA VIA12_2cut_HN DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M1 ;
        RECT -0.050 -0.090  0.050  0.330 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.190  0.050  0.290 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.330 ;
END VIA12_2cut_HN

VIA VIA12_2cut_HS DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M1 ;
        RECT -0.050 -0.330  0.050  0.090 ;
    LAYER VIA1 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.290  0.050 -0.190 ;
    LAYER M2 ;
        RECT -0.050 -0.330  0.050  0.090 ;
END VIA12_2cut_HS

VIA VIA12_4cut DEFAULT
    RESISTANCE 0.3750000000 ;
    LAYER M1 ;
        RECT -0.190 -0.150  0.190  0.150 ;
    LAYER VIA1 ;
        RECT -0.150 -0.150 -0.050 -0.050 ;
        RECT -0.150  0.050 -0.050  0.150 ;
        RECT  0.050  0.050  0.150  0.150 ;
        RECT  0.050 -0.150  0.150 -0.050 ;
    LAYER M2 ;
        RECT -0.150 -0.190  0.150  0.190 ;
END VIA12_4cut

VIA VIA23_1cut DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA23_1cut

VIA VIA23_1cut_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA23_1cut_V
                 
VIA VIA23_1cut_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA23_1cut_H

VIA VIA23_1cut_FAT_C DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA23_1cut_FAT_C
             
VIA VIA23_1cut_FAT_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA23_1cut_FAT_V

VIA VIA23_1cut_FAT_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA23_1cut_FAT_H

VIA VIA23_1cut_FAT DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.090 -0.090  0.090  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.090  0.090  0.090 ;
END VIA23_1cut_FAT
                 
VIA VIA23_1stack_N DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.430 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA23_1stack_N

VIA VIA23_1stack_S DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M2 ;
        RECT -0.050 -0.430  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA23_1stack_S

VIA VIA23_2cut_E DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.250  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.290  0.050 ;
END VIA23_2cut_E

VIA VIA23_2cut_W DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M2 ;
        RECT -0.250 -0.090  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M3 ;
        RECT -0.290 -0.050  0.090  0.050 ;
END VIA23_2cut_W

VIA VIA23_2cut_N DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M2 ;
        RECT -0.050 -0.090  0.050  0.290 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.250 ;
END VIA23_2cut_N

VIA VIA23_2cut_S DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M2 ;
        RECT -0.050 -0.290  0.050  0.090 ;
    LAYER VIA2 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M3 ;
        RECT -0.090 -0.250  0.090  0.050 ;
END VIA23_2cut_S

VIA VIA23_4cut DEFAULT
    RESISTANCE 0.3750000000 ;
    LAYER M2 ;
        RECT -0.150 -0.190  0.150  0.190 ;
    LAYER VIA2 ;
        RECT -0.150 -0.150 -0.050 -0.050 ;
        RECT -0.150  0.050 -0.050  0.150 ;
        RECT  0.050  0.050  0.150  0.150 ;
        RECT  0.050 -0.150  0.150 -0.050 ;
    LAYER M3 ;
        RECT -0.190 -0.150  0.190  0.150 ;
END VIA23_4cut

VIA VIA34_1cut DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA34_1cut

VIA VIA34_1cut_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA34_1cut_H
                 
VIA VIA34_1cut_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA34_1cut_V

VIA VIA34_1cut_FAT_C DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA34_1cut_FAT_C
             
VIA VIA34_1cut_FAT_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA34_1cut_FAT_H

VIA VIA34_1cut_FAT_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA34_1cut_FAT_V

VIA VIA34_1cut_FAT DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.090 -0.090  0.090  0.090 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.090 -0.090  0.090  0.090 ;
END VIA34_1cut_FAT
                 
VIA VIA34_1stack_E DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.430  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA34_1stack_E

VIA VIA34_1stack_W DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M3 ;
        RECT -0.430 -0.050  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA34_1stack_W

VIA VIA34_2cut_E DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.290  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.250  0.090 ;
END VIA34_2cut_E

VIA VIA34_2cut_W DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M3 ;
        RECT -0.290 -0.050  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M4 ;
        RECT -0.250 -0.090  0.050  0.090 ;
END VIA34_2cut_W

VIA VIA34_2cut_N DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M3 ;
        RECT -0.090 -0.050  0.090  0.250 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.290 ;
END VIA34_2cut_N

VIA VIA34_2cut_S DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M3 ;
        RECT -0.090 -0.250  0.090  0.050 ;
    LAYER VIA3 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M4 ;
        RECT -0.050 -0.290  0.050  0.090 ;
END VIA34_2cut_S

VIA VIA34_4cut DEFAULT
    RESISTANCE 0.3750000000 ;
    LAYER M3 ;
        RECT -0.190 -0.150  0.190  0.150 ;
    LAYER VIA3 ;
        RECT -0.150 -0.150 -0.050 -0.050 ;
        RECT -0.150  0.050 -0.050  0.150 ;
        RECT  0.050  0.050  0.150  0.150 ;
        RECT  0.050 -0.150  0.150 -0.050 ;
    LAYER M4 ;
        RECT -0.150 -0.190  0.150  0.190 ;
END VIA34_4cut

VIA VIA45_1cut DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA45_1cut

VIA VIA45_1cut_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA45_1cut_V
                 
VIA VIA45_1cut_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA45_1cut_H

VIA VIA45_1cut_FAT_C DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA45_1cut_FAT_C
             
VIA VIA45_1cut_FAT_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA45_1cut_FAT_V

VIA VIA45_1cut_FAT_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA45_1cut_FAT_H

VIA VIA45_1cut_FAT DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.090 -0.090  0.090  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.090  0.090  0.090 ;
END VIA45_1cut_FAT
                 
VIA VIA45_1stack_N DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.430 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA45_1stack_N

VIA VIA45_1stack_S DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M4 ;
        RECT -0.050 -0.430  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA45_1stack_S

VIA VIA45_2cut_E DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.250  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.290  0.050 ;
END VIA45_2cut_E

VIA VIA45_2cut_W DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M4 ;
        RECT -0.250 -0.090  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M5 ;
        RECT -0.290 -0.050  0.090  0.050 ;
END VIA45_2cut_W

VIA VIA45_2cut_N DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M4 ;
        RECT -0.050 -0.090  0.050  0.290 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.250 ;
END VIA45_2cut_N

VIA VIA45_2cut_S DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M4 ;
        RECT -0.050 -0.290  0.050  0.090 ;
    LAYER VIA4 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M5 ;
        RECT -0.090 -0.250  0.090  0.050 ;
END VIA45_2cut_S

VIA VIA45_4cut DEFAULT
    RESISTANCE 0.3750000000 ;
    LAYER M4 ;
        RECT -0.150 -0.190  0.150  0.190 ;
    LAYER VIA4 ;
        RECT -0.150 -0.150 -0.050 -0.050 ;
        RECT -0.150  0.050 -0.050  0.150 ;
        RECT  0.050  0.050  0.150  0.150 ;
        RECT  0.050 -0.150  0.150 -0.050 ;
    LAYER M5 ;
        RECT -0.190 -0.150  0.190  0.150 ;
END VIA45_4cut

VIA VIA56_1cut DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA56_1cut

VIA VIA56_1cut_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.090 -0.050  0.090  0.050 ;
END VIA56_1cut_H
                 
VIA VIA56_1cut_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.050 -0.090  0.050  0.090 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA56_1cut_V

VIA VIA56_1cut_FAT_C DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA56_1cut_FAT_C
             
VIA VIA56_1cut_FAT_H DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.12 -0.050  0.12  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.12 -0.050  0.12  0.050 ;
END VIA56_1cut_FAT_H

VIA VIA56_1cut_FAT_V DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.050 -0.12  0.050  0.12 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.12  0.050  0.12 ;
END VIA56_1cut_FAT_V

VIA VIA56_1cut_FAT DEFAULT
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.090 -0.090  0.090  0.090 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.090 -0.090  0.090  0.090 ;
END VIA56_1cut_FAT
                 
VIA VIA56_1stack_E DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.430  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA56_1stack_E

VIA VIA56_1stack_W DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.5000000000 ;
    LAYER M5 ;
        RECT -0.430 -0.050  0.090  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.090  0.050  0.090 ;
END VIA56_1stack_W

VIA VIA56_2cut_E DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.290  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.090  0.250  0.090 ;
END VIA56_2cut_E

VIA VIA56_2cut_W DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M5 ;
        RECT -0.290 -0.050  0.090  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M6 ;
        RECT -0.250 -0.090  0.050  0.090 ;
END VIA56_2cut_W

VIA VIA56_2cut_N DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.090  0.250 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050  0.150  0.050  0.250 ;
    LAYER M6 ;
        RECT -0.050 -0.090  0.050  0.290 ;
END VIA56_2cut_N

VIA VIA56_2cut_S DEFAULT
    RESISTANCE 0.7500000000 ;
    LAYER M5 ;
        RECT -0.090 -0.250  0.090  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.050 -0.250  0.050 -0.150 ;
    LAYER M6 ;
        RECT -0.050 -0.290  0.050  0.090 ;
END VIA56_2cut_S

VIA VIA56_2stack_E DEFAULT TOPOFSTACKONLY
    RESISTANCE 0.7500000000 ;
    LAYER M5 ;
        RECT -0.090 -0.050  0.430  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT  0.150 -0.050  0.250  0.050 ;
    LAYER M6 ;
        RECT -0.050 -0.090  0.250  0.090 ;
END VIA56_2stack_E
 
VIA VIA56_2stack_W DEFAULT TOPOFSTACKONLY
    RESISTANCE 0.7500000000 ;
    LAYER M5 ;
        RECT -0.430 -0.050  0.090  0.050 ;
    LAYER VIA5 ;
        RECT -0.050 -0.050  0.050  0.050 ;
        RECT -0.250 -0.050 -0.150  0.050 ;
    LAYER M6 ;
        RECT -0.250 -0.090  0.050  0.090 ;
END VIA56_2stack_W

VIA VIA56_4cut DEFAULT
    RESISTANCE 0.3750000000 ;
    LAYER M5 ;
        RECT -0.190 -0.150  0.190  0.150 ;
    LAYER VIA5 ;
        RECT -0.150 -0.150 -0.050 -0.050 ;
        RECT -0.150  0.050 -0.050  0.150 ;
        RECT  0.050  0.050  0.150  0.150 ;
        RECT  0.050 -0.150  0.150 -0.050 ;
    LAYER M6 ;
        RECT -0.150 -0.190  0.150  0.190 ;
END VIA56_4cut

VIA VIA67_1cut DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.200  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
END VIA67_1cut
 
VIA VIA67_1cut_V DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.200  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA67_1cut_V
 
VIA VIA67_1cut_H DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M6 ;
        RECT -0.260 -0.200  0.260  0.200 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
END VIA67_1cut_H
 
VIA VIA67_1cut_FAT_C DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M6 ;
        RECT -0.200 -0.26  0.200  0.26 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.26 -0.200  0.26  0.200 ;
END VIA67_1cut_FAT_C
 
VIA VIA67_1cut_FAT_V DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M6 ;
        RECT -0.200 -0.26  0.200  0.26 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.200 -0.26  0.200  0.26 ;
END VIA67_1cut_FAT_V
 
VIA VIA67_1cut_FAT_H DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M6 ;
        RECT -0.26 -0.200  0.26  0.200 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.26 -0.200  0.26  0.200 ;
END VIA67_1cut_FAT_H
 
VIA VIA67_1cut_FAT DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M6 ;
        RECT -0.260 -0.260  0.260  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M7 ;
        RECT -0.260 -0.260  0.260  0.260 ;
END VIA67_1cut_FAT
 
VIA VIA67_2cut_E DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.900  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT  0.520 -0.180  0.880  0.180 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.960  0.200 ;
END VIA67_2cut_E
 
VIA VIA67_2cut_W DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M6 ;
        RECT -0.900 -0.260  0.200  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.880 -0.180 -0.520  0.180 ;
    LAYER M7 ;
        RECT -0.960 -0.200  0.260  0.200 ;
END VIA67_2cut_W
 
VIA VIA67_2cut_N DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M6 ;
        RECT -0.200 -0.260  0.200  0.960 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.180  0.520  0.180  0.880 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.900 ;
END VIA67_2cut_N
 
VIA VIA67_2cut_S DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M6 ;
        RECT -0.200 -0.960  0.200  0.260 ;
    LAYER VIA6 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.180 -0.880  0.180 -0.520 ;
    LAYER M7 ;
        RECT -0.260 -0.900  0.260  0.200 ;
END VIA67_2cut_S
 
VIA VIA67_4cut DEFAULT
    RESISTANCE 0.0550000000 ;
    LAYER M6 ;
        RECT -0.650 -0.710  0.650  0.710 ;
    LAYER VIA6 ;
        RECT -0.630 -0.630 -0.270 -0.270 ;
        RECT -0.630  0.270 -0.270  0.630 ;
        RECT  0.270  0.270  0.630  0.630 ;
        RECT  0.270 -0.630  0.630 -0.270 ;
    LAYER M7 ;
        RECT -0.710 -0.650  0.710  0.650 ;
END VIA67_4cut

VIA VIA78_1cut DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA78_1cut
 
VIA VIA78_1cut_H DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.260 -0.200  0.260  0.200 ;
END VIA78_1cut_H
 
VIA VIA78_1cut_V DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.200 -0.260  0.200  0.260 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA78_1cut_V
 
VIA VIA78_1cut_FAT_C DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.26 -0.200  0.26  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.26  0.200  0.26 ;
END VIA78_1cut_FAT_C
 
VIA VIA78_1cut_FAT_H DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.26 -0.200  0.26  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.26 -0.200  0.26  0.200 ;
END VIA78_1cut_FAT_H
 
VIA VIA78_1cut_FAT_V DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.200 -0.26  0.200  0.26 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.26  0.200  0.26 ;
END VIA78_1cut_FAT_V
 
VIA VIA78_1cut_FAT DEFAULT
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.260 -0.260  0.260  0.260 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.260 -0.260  0.260  0.260 ;
END VIA78_1cut_FAT

VIA VIA78_1stack_E DEFAULT TOPOFSTACKONLY
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  1.155  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA78_1stack_E
 
VIA VIA78_1stack_W DEFAULT TOPOFSTACKONLY
    RESISTANCE 0.2200000000 ;
    LAYER M7 ;
        RECT -1.155 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.260 ;
END VIA78_1stack_W
 
VIA VIA78_2cut_E DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.960  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT  0.520 -0.180  0.880  0.180 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.900  0.260 ;
END VIA78_2cut_E
 
VIA VIA78_2cut_W DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M7 ;
        RECT -0.960 -0.200  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.880 -0.180 -0.520  0.180 ;
    LAYER M8 ;
        RECT -0.900 -0.260  0.200  0.260 ;
END VIA78_2cut_W
 
VIA VIA78_2cut_N DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M7 ;
        RECT -0.260 -0.200  0.260  0.900 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.180  0.520  0.180  0.880 ;
    LAYER M8 ;
        RECT -0.200 -0.260  0.200  0.960 ;
END VIA78_2cut_N
 
VIA VIA78_2cut_S DEFAULT
    RESISTANCE 0.1100000000 ;
    LAYER M7 ;
        RECT -0.260 -0.900  0.260  0.200 ;
    LAYER VIA7 ;
        RECT -0.180 -0.180  0.180  0.180 ;
        RECT -0.180 -0.880  0.180 -0.520 ;
    LAYER M8 ;
        RECT -0.200 -0.960  0.200  0.260 ;
END VIA78_2cut_S
 
VIA VIA78_4cut DEFAULT
    RESISTANCE 0.0550000000 ;
    LAYER M7 ;
        RECT -0.710 -0.650  0.710  0.650 ;
    LAYER VIA7 ;
        RECT -0.630 -0.630 -0.270 -0.270 ;
        RECT -0.630  0.270 -0.270  0.630 ;
        RECT  0.270  0.270  0.630  0.630 ;
        RECT  0.270 -0.630  0.630 -0.270 ;
    LAYER M8 ;
        RECT -0.650 -0.710  0.650  0.710 ;
END VIA78_4cut
 
VIARULE VIAGEN12 GENERATE
    LAYER M1 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.09 TO 12.00 ;
    LAYER M2 ;
        ENCLOSURE 0.4E-01 0 ;
        WIDTH 0.10 TO 12.00 ;
    LAYER VIA1 ;
        RECT -0.5E-01 -0.5E-01 0.5E-01 0.5E-01 ;
        SPACING 0.23 BY 0.23 ;    
END VIAGEN12        

VIARULE VIAGEN23 GENERATE
    LAYER M2 ;
        ENCLOSURE 0.4E-01 0 ;  
        WIDTH 0.10 TO 12.00 ;
    LAYER M3 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER VIA2 ;
        RECT -0.5E-01 -0.5E-01 0.5E-01 0.5E-01 ; 
        SPACING 0.23 BY 0.23 ;    
END VIAGEN23

VIARULE VIAGEN34 GENERATE
    LAYER M3 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER M4 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER VIA3 ;
        RECT -0.5E-01 -0.5E-01 0.5E-01 0.5E-01 ; 
        SPACING 0.23 BY 0.23 ;    
END VIAGEN34

VIARULE VIAGEN45 GENERATE
    LAYER M4 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER M5 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER VIA4 ;
        RECT -0.5E-01 -0.5E-01 0.5E-01 0.5E-01 ; 
        SPACING 0.23 BY 0.23 ;    
END VIAGEN45

VIARULE VIAGEN56 GENERATE
    LAYER M5 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER M6 ;
        ENCLOSURE 0.4E-01 0 ; 
        WIDTH 0.10 TO 12.00 ;
    LAYER VIA5 ;
        RECT -0.5E-01 -0.5E-01 0.5E-01 0.5E-01 ; 
        SPACING 0.23 BY 0.23 ;    
END VIAGEN56

VIARULE VIAGEN67 GENERATE
    LAYER M6 ;
        ENCLOSURE 0.8E-01 0.2E-01  ;
        WIDTH 0.10 TO 12.00 ;
    LAYER M7 ;
        ENCLOSURE 0.8E-01 0.2E-01  ;
        WIDTH 0.40 TO 12.00 ;
    LAYER VIA6 ;
        RECT -0.18 -0.18 0.18 0.18 ; 
        SPACING 0.90 BY 0.90 ;    
END VIAGEN67

VIARULE VIAGEN78 GENERATE
    LAYER M7 ;
        ENCLOSURE 0.8E-01 0.2E-01  ;
        WIDTH 0.40 TO 12.00 ;
    LAYER M8 ;
        ENCLOSURE 0.8E-01 0.2E-01  ;
        WIDTH 0.40 TO 12.00 ;
    LAYER VIA7 ;
        RECT -0.18 -0.18 0.18 0.18 ; 
        SPACING 0.90 BY 0.90 ;    
END VIAGEN78           

MAXVIASTACK 4 RANGE M1 M6 ;

VIARULE TURN1 GENERATE
    LAYER M1 ;
        DIRECTION HORIZONTAL ;
    LAYER M1 ;
        DIRECTION VERTICAL ;
END TURN1

VIARULE TURN2 GENERATE
    LAYER M2 ;
        DIRECTION HORIZONTAL ;
    LAYER M2 ;
        DIRECTION VERTICAL ;
END TURN2

VIARULE TURN3 GENERATE
    LAYER M3 ;
        DIRECTION HORIZONTAL ;
    LAYER M3 ;
        DIRECTION VERTICAL ;
END TURN3

VIARULE TURN4 GENERATE
    LAYER M4 ;
        DIRECTION HORIZONTAL ;
    LAYER M4 ;
        DIRECTION VERTICAL ;
END TURN4

VIARULE TURN5 GENERATE
    LAYER M5 ;
        DIRECTION HORIZONTAL ;
    LAYER M5 ;
        DIRECTION VERTICAL ;
END TURN5

VIARULE TURN6 GENERATE
    LAYER M6 ;
        DIRECTION HORIZONTAL ;
    LAYER M6 ;
        DIRECTION VERTICAL ;
END TURN6

VIARULE TURN7 GENERATE
    LAYER M7 ;
        DIRECTION HORIZONTAL ;
    LAYER M7 ;
        DIRECTION VERTICAL ;
END TURN7

VIARULE TURN8 GENERATE
    LAYER M8 ;
        DIRECTION HORIZONTAL ;
    LAYER M8 ;
        DIRECTION VERTICAL ;
END TURN8

SITE core
    SIZE 0.20 BY 1.80 ;
    CLASS CORE ;
    SYMMETRY Y  ;
END core

SITE bcore
    SIZE 0.20 BY 3.60 ;
    CLASS CORE ;
    SYMMETRY Y  ;
END bcore
 
SITE ccore
    SIZE 0.20 BY 5.40 ;
    CLASS CORE ;
    SYMMETRY Y  ;
END ccore
 
SITE dcore
    SIZE 0.20 BY 7.20 ;
    CLASS CORE ;
    SYMMETRY Y  ;
END dcore
 
SITE gacore
    SIZE 0.80 BY 1.80 ;
    CLASS CORE ;
    SYMMETRY Y  ;
END gacore

END LIBRARY
